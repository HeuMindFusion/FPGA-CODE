module multiply (y,a,b);
input [7:0] a,b;
ouput reg [7:0] y;
always @(a or b)
begin
y[0]<=(a[0]&a[0])^(a[1]&a[7])^(a[2]&a[6])^(a[3]&a[5])^(a[4]&a[4])^(a[5]&a[3])^(a[6]&a[2])^(a[7]&a[1])^
	       (a[5]&a[7])^(a[6]&a[6])^(a[7]&a[5])^(a[6]&a[7])^(a[7]&a[6])^(a[7]&a[7]);	
	 y[1]<=(a[0]&a[1])^(a[1]&a[0])^(a[2]&a[7])^(a[3]&a[6])^(a[4]&a[5])^(a[5]&a[4])^(a[6]&a[3])^(a[7]&a[2])^
	      (a[6]&a[7])^(a[7]&a[6])^(a[7]&a[7]);	
y[2]<=(a[0]&a[2])^(a[1]&a[1])^(a[2]&a[0])^(a[1]&a[7])^(a[2]&a[6])^(a[3]&a[5])^(a[4]&a[4])^(a[5]&a[3])^
	       (a[6]&a[2])^(a[7]&a[1])^(a[3]&a[7])^(a[4]&a[6])^(a[5]&a[5])^(a[6]&a[4])^(a[7]&a[3])^(a[5]&a[7])^
	       (a[6]&a[6])^(a[7]&a[5])^(a[6]&a[7])^(a[7]&a[6]);	
      y[3]<=(a[0]&a[3])^(a[1]&a[2])^(a[2]&a[1])^(a[3]&a[0])^(a[1]&a[7])^(a[2]&a[6])^(a[3]&a[5])^(a[4]&a[4])^
	       (a[5]&a[3])^(a[6]&a[2])^(a[7]&a[1])^(a[2]&a[7])^(a[3]&a[6])^(a[4]&a[5])^(a[5]&a[4])^(a[6]&a[3])^
		  (a[7]&a[2])^(a[4]&a[7])^(a[5]&a[6])^(a[6]&a[5])^(a[7]&a[4])^(a[5]&a[7])^(a[6]&a[6])^(a[7]&a[5]);	
    y[4]<=(a[0]&a[4])^(a[1]&a[3])^(a[2]&a[2])^(a[3]&a[1])^(a[4]&a[0])^(a[1]&a[7])^(a[2]&a[6])^(a[3]&a[5])^
	     (a[4]&a[4])^(a[5]&a[3])^(a[6]&a[2])^(a[7]&a[1])^(a[2]&a[7])^(a[3]&a[6])^(a[4]&a[5])^(a[5]&a[4])^
	     (a[6]&a[3])^(a[7]&a[2])^(a[3]&a[7])^(a[4]&a[6])^(a[5]&a[5])^(a[6]&a[4])^(a[7]&a[3])^(a[7]&a[7]);	
	 y[5]<=(a[0]&a[5])^(a[1]&a[4])^(a[2]&a[3])^(a[3]&a[2])^(a[4]&a[1])^(a[5]&a[0])^(a[2]&a[7])^(a[3]&a[6])^
	      (a[4]&a[5])^(a[5]&a[4])^(a[6]&a[3])^(a[7]&a[2])^(a[3]&a[7])^(a[4]&a[6])^(a[5]&a[5])^(a[6]&a[4])^
		  (a[7]&a[3])^(a[4]&a[7])^(a[5]&a[6])^(a[6]&a[5])^(a[7]&a[4]);	
	 y[6]<=(a[0]&a[6])^(a[1]&a[5])^(a[2]&a[4])^(a[3]&a[3])^(a[4]&a[2])^(a[5]&a[1])^(a[6]&a[0])^(a[3]&a[7])^
	       (a[4]&a[6])^(a[5]&a[5])^(a[6]&a[4])^(a[7]&a[3])^(a[4]&a[7])^(a[5]&a[6])^(a[6]&a[5])^(a[7]&a[4])^
		  (a[5]&a[7])^(a[6]&a[6])^(a[7]&a[5]);	
	 y[7]<=(a[0]&a[7])^(a[1]&a[6])^(a[2]&a[5])^(a[3]&a[4])^(a[4]&a[3])^(a[5]&a[2])^(a[6]&a[1])^(a[7]&a[0])^
	       (a[4]&a[7])^(a[5]&a[6])^(a[6]&a[5])^(a[7]&a[4])^(a[7]&a[6])^(a[5]&a[7])^(a[6]&a[6])^(a[7]&a[5])^
		  (a[6]&a[7])^(a[7]&a[6]);
end
endmodule
