`timescale 1ns / 1ps


module ldpc(clk,data,out);
input clk;
input data;
output reg out;
//A
reg [10:0] addra=11'd0;
wire [8:0] douta;
//C
reg[6:0]addra1=7'd0;
wire[8:0]douta1;
//ETT
reg[8:0]addra2=9'd0;
wire[8:0]douta2;
//p
reg[5:0]addra3=6'd0;
wire[4:0]douta3;
//TT
reg[10:0]addra4=11'd0;
wire[8:0]douta4;

reg [263:0]au;
reg [23:0]cu;
reg [23:0]tu;
reg [23:0]p1;
reg [263:0]bp1;
reg [263:0]bp2;
reg [263:0]p2;

reg[287:0]u;//������Ϣλ
reg[575:0]u1;//��������
reg [4:0]a;
reg [3:0]b;
reg[10:0]c;
reg[10:0]d;

reg[8:0]j=9'd0;//au����������
reg[8:0]cnt=9'd0;//������Ϣ����ȼ��?reg[2:0]i=3'd0;//����a��u��Ӧ1��λ�õļ�����
reg[3:0]i1=4'd0;//����c��au��Ӧ1��λ�õļ�����

reg [7:0]k=8'd0;//����λ��

reg[4:0]j1=5'd0;//cu���м�����
reg[4:0]j2=5'd0;//et��au���м�����
reg[8:0]j3=9'd0;
reg[9:0]j4=10'd0;

reg[4:0]i2=5'd0;//et��au����cuʱ��λ������
reg[8:0]i3=9'd0;
reg[8:0]i4=9'd0;
reg[3:0]i5=4'd0;

A  a1_2(.clka(clk),.addra(addra),.douta(douta));
C  c1_2(.clka(clk),.addra(addra1),.douta(douta1));
ETT ett1_2(.clka(clk),.addra(addra2),.douta(douta2));
p  p1_2(.clka(clk),.addra(addra3),.douta(douta3));
TT tt1_2(.clka(clk),.addra(addra4),.douta(douta4));

//k1=k30 result au
always@(posedge clk)
case(k)
 8'd0:begin//��ʼ��������Ϣλu
  if(cnt<9'd288)
  begin
   cnt<=cnt+1; 
  u<={data,u[287:1]};
  end
  else
  k<=8'd1;
  end
 8'd1:begin
   a[i]<=u[douta];
	b[i]<=u[douta1];
	k<=8'd2;
	end	
 8'd2:begin  
   addra<=addra+1;
	addra1<=addra1+1;
	k<=8'd3;
	end
 8'd3:begin 
    if(i<3)
	 begin 
	  i<=i+1;
	  k<=8'd1;
	  end
	  else
	  k<=8'd4;
	  end	  
  8'd4:begin 
   au[j]<=a[0]^a[1]^a[2]^a[3];
	cu[j1]<=b[0]^b[1]^b[2]^b[3];
	k<=8'd5;
	end	
	8'd5:begin 
	    j<=j+1;
		 j1<=j1+1;
		 i<=3'd0;
		 k<=8'd6;
		 end		 
	 8'd6:begin 
       if(j<=9'd23) 
	    k<=8'd1;
	    else
	     k<=8'd7;
	     end	  
	 8'd7:begin
        a[i]<=u[douta];
	     k<=8'd8;
	      end	
   8'd8:begin  
        addra<=addra+1;
	      k<=8'd9;
	     end
   8'd9:begin 
        if(i<4)
	      begin 
	      i<=i+1;
	      k<=8'd7;
	      end
	      else
	      k<=8'd10;
	      end	  
    8'd10:begin 
         au[j]<=a[0]^a[1]^a[2]^a[3]^a[4];
	      k<=8'd11;
	       end	
	  8'd11:begin 
	    j<=j+1;
		 i<=3'd0;
		 k<=8'd12;
		 end	 
	  8'd12:begin 
       if(j<=9'd71) 
	    k<=8'd7;
	   else
	   begin
	   k<=8'd13;
	   end
	   end		
   8'd13:begin
      a[i]<=u[douta];
	   k<=8'd14;
	   end
   8'd14:begin  
        addra<=addra+1;
	     k<=8'd15;
	     end
   8'd15:begin 
        if(i<3)
	     begin 
	     i<=i+1;
	     k<=8'd13;
	     end
	     else
	     k<=8'd16;
	     end  
    8'd16:begin 
       au[j]<=a[0]^a[1]^a[2]^a[3];
	    k<=8'd17;
	    end
	 8'd17:begin 
	    j<=j+1;
		 i<=3'd0;
		 k<=8'd18;
		 end	 
	 8'd18:begin 
       if(j<=9'd191) 
	    k<=8'd13;
	    else
	    k<=8'd19;
	    end		  
	 8'd19:begin
        a[i]<=u[douta];
	     k<=8'd20;
	      end	
   8'd20:begin  
        addra<=addra+1;
	      k<=8'd21;
	     end
   8'd21:begin 
        if(i<4)
	      begin 
	      i<=i+1;
	      k<=8'd19;
	      end
	      else
	      k<=8'd22;
	      end	  
    8'd22:begin 
         au[j]<=a[0]^a[1]^a[2]^a[3]^a[4];
	      k<=8'd23;
	       end	
	  8'd23:begin 
	    j<=j+1;
		 i<=3'd0;
		 k<=8'd24;
		 end		 
	  8'd24:begin 
       if(j<=9'd215) 
	    k<=8'd19;
	   else
	   begin
	   k<=8'd25;
	   end
	   end		
		8'd25:begin
        a[i]<=u[douta];
	     k<=8'd26;
	     end	
     8'd26:begin  
         addra<=addra+1;
	      k<=8'd27;
	      end
     8'd27:begin 
        if(i<3)
	     begin 
	     i<=i+1;
	     k<=8'd25;
	     end
	     else
	     k<=8'd28;
	     end	  
     8'd28:begin 
        au[j]<=a[0]^a[1]^a[2]^a[3];
	     k<=8'd29;
	     end	
	  8'd29:begin 
	    j<=j+1;
		 i<=3'd0;
		 k<=8'd30;
		 end		 
	  8'd30:begin 
       if(j<=9'd263) 
	    k<=8'd25;
	    else
	     k<=8'd31;
	     end
	//p1	  	
   8'd31:begin
      c[i1]<=au[douta2];
	   k<=8'd32;
	   end	
   8'd32:begin  
        addra2<=addra2+1;
	     k<=8'd33;
	     end
   8'd33:begin 
        if(i1<10)
	     begin 
	     i1<=i1+1;
	     k<=8'd31;
	     end
	     else
	     k<=8'd34;
	     end	  
    8'd34:begin 
       tu[j2]<=c[0]^c[1]^c[2]^c[3]^c[4]^c[5]^c[6]^c[7]^c[8]^c[9]^c[10];
	    k<=8'd35;
	    end	
	 8'd35:begin 
	    j2<=j2+1;
		 i1<=4'd0;
		 k<=8'd36;
		 end	 
	 8'd36:begin 
       if(j2<=5'd23) 
	    k<=8'd31;
	    else
	    k<=8'd37;
	    end
	 8'd37:begin
			 p1[i2]<=tu[i2]^cu[i2];
			  k<=8'd38;
				end
	 8'd38:begin 
	        if(i2<23)
			  begin 
			   i2<=i2+1;
				k<=8'd37;
				end
				else
				k<=8'd39;
				end
	//B*p1
	  8'd39:begin
			 if(i3<24||(119<i3&&i3<144))//У�����1������λ��
			 begin 
			 bp1[i3]<=p1[douta3];
			 k<=8'd40;
			 end
			 else
			 begin 
			 bp1[i3]<=0;
			 k<=8'd41;
			 end
			 end
		8'd40:begin 
		      addra3<=addra3+1;
				k<=8'd41;
				end
		8'd41:begin 
		      if(i3<264)
				  begin 
				  i3<=i3+1;
				  k<=8'd39;
				  end
				 else
				   k<=8'd42;
					end
	//au+bp1;
	    8'd42:begin
			 bp2[i4]<=bp1[i4]^au[i4];
			  k<=8'd43;
				end
	    8'd43:begin 
	        if(i4<263)
			  begin 
			   i4<=i4+1;
				k<=8'd42;
				end
				else
				k<=8'd44;
				end
		//p2
	   8'd44:begin//��һ��
        p2[j3]<=bp2[douta4];
	     k<=8'd45;
	      end
      8'd45:begin  
        addra4<=addra4+1;
	      k<=8'd46;
	     end
       8'd46:begin 
        if(j3<23)
	      begin 
	      j3<=j3+1;
	      k<=8'd44;
	      end
	      else
			begin
			j3<=j3+1;
	      k<=8'd47;
			end
	      end		
		8'd47:begin//�ڶ��п�ʼ
        d[i5]<=bp2[douta4];
	     k<=8'd48;
	      end
      8'd48:begin  
        addra4<=addra4+1;
	      k<=8'd49;
	     end
      8'd49:begin 
        if(i5<1)
	      begin 
	      i5<=i5+1;
	      k<=8'd47;
	      end
	      else
	      k<=8'd50;
	      end 
      8'd50:begin 
         p2[j3]<=d[0]^d[1];
	      k<=8'd51;
	       end
	   8'd51:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd52;
		 end	 
      8'd52:begin 
       if(j3<=9'd47) //////////////////////////////////
	    k<=8'd47;
	   else
	   begin
	   k<=8'd53;
	   end
	   end	
      8'd53:begin
        d[i5]<=bp2[douta4];
	     k<=8'd54;
	      end
      8'd54:begin  
        addra4<=addra4+1;
	      k<=8'd55;
	     end
      8'd55:begin 
        if(i5<2)
	      begin 
	      i5<=i5+1;
	      k<=8'd53;
	      end
	      else
	      k<=8'd56;
	      end  
      8'd56:begin 
         p2[j3]<=d[0]^d[1]^d[2];
	      k<=8'd57;
	       end
	   8'd57:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd58;
		 end	 
	   8'd58:begin 
       if(j3<=9'd71) 
	    k<=8'd53;
	   else
	   begin
	   k<=8'd59;
	   end
	   end	
      8'd59:begin
        d[i5]<=bp2[douta4];
	     k<=8'd60;
	      end
      8'd60:begin  
        addra4<=addra4+1;
	      k<=8'd61;
	     end
      8'd61:begin 
        if(i5<3)
	      begin 
	      i5<=i5+1;
	      k<=8'd59;
	      end
	      else
	      k<=8'd62;
	      end 
      8'd62:begin 
         p2[j3]<=d[0]^d[1]^d[2]^d[3];
	      k<=8'd63;
	       end
	   8'd63:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd64;
		 end 
	   8'd64:begin 
       if(j3<=9'd95) 
	    k<=8'd59;
	   else
	   begin
	   k<=8'd65;
	   end
	   end	
      8'd65:begin
        d[i5]<=bp2[douta4];
	     k<=8'd66;
	      end
      8'd66:begin  
        addra4<=addra4+1;
	      k<=8'd67;
	     end
      8'd67:begin 
        if(i5<4)
	      begin 
	      i5<=i5+1;
	      k<=8'd65;
	      end
	      else
	      k<=8'd68;
	      end 
      8'd68:begin 
         p2[j3]<=d[0]^d[1]^d[2]^d[3]^d[4];
	      k<=8'd69;
	       end
	   8'd69:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd70;
		 end		 
	   8'd70:begin 
       if(j3<=9'd119) 
	    k<=8'd65;
	   else
	   begin
	   k<=8'd71;
	   end
	   end
		 8'd71:begin
        d[i5]<=bp2[douta4];
	     k<=8'd72;
	      end
      8'd72:begin  
        addra4<=addra4+1;
	      k<=8'd73;
	     end
      8'd73:begin 
        if(i5<5)
	      begin 
	      i5<=i5+1;
	      k<=8'd71;
	      end
	      else
	      k<=8'd74;
	      end	  
      8'd74:begin 
         p2[j3]<=d[0]^d[1]^d[2]^d[3]^d[4]^d[5];
	      k<=8'd75;
	       end
	   8'd75:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd76;
		 end	 
	   8'd76:begin 
       if(j3<=9'd143) 
	    k<=8'd71;
	   else
	   begin
	   k<=8'd77;
	   end
	   end	
		 8'd77:begin
        d[i5]<=bp2[douta4];
	     k<=8'd78;
	      end
      8'd78:begin  
        addra4<=addra4+1;
	      k<=8'd79;
	     end
      8'd79:begin 
        if(i5<6)
	      begin 
	      i5<=i5+1;
	      k<=8'd77;
	      end
	      else
	      k<=8'd80;
	      end  
      8'd80:begin 
         p2[j3]<=d[0]^d[1]^d[2]^d[3]^d[4]^d[5]^d[6];
	      k<=8'd81;
	       end
	   8'd81:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd82;
		 end	 
	   8'd82:begin 
       if(j3<=9'd167) 
	    k<=8'd77;
	   else
	   begin
	   k<=8'd83;
	   end
	   end	
		 8'd83:begin
        d[i5]<=bp2[douta4];
	     k<=8'd84;
	      end
      8'd84:begin  
        addra4<=addra4+1;
	      k<=8'd85;
	     end
      8'd85:begin 
        if(i5<7)
	      begin 
	      i5<=i5+1;
	      k<=8'd83;
	      end
	      else
	      k<=8'd86;
	      end 
      8'd86:begin 
         p2[j3]<=d[0]^d[1]^d[2]^d[3]^d[4]^d[5]^d[6]^d[7];
	      k<=8'd87;
	       end
	   8'd87:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd88;
		 end		 
	   8'd88:begin 
       if(j3<=9'd191) 
	    k<=8'd83;
	   else
	   begin
	   k<=8'd89;
	   end
	   end	
		8'd89:begin
        d[i5]<=bp2[douta4];
	     k<=8'd90;
	      end
      8'd90:begin  
        addra4<=addra4+1;
	      k<=8'd91;
	     end
      8'd91:begin 
        if(i5<8)
	      begin 
	      i5<=i5+1;
	      k<=8'd89;
	      end
	      else
	      k<=8'd92;
	      end
      8'd92:begin 
         p2[j3]<=d[0]^d[1]^d[2]^d[3]^d[4]^d[5]^d[6]^d[7]^d[8];
	      k<=8'd93;
	       end
	   8'd93:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd94;
		 end	 
	   8'd94:begin 
       if(j3<=9'd215) 
	    k<=8'd89;
	   else
	   begin
	   k<=8'd95;
	   end
	   end
		8'd95:begin
        d[i5]<=bp2[douta4];
	     k<=8'd96;
	      end
      8'd96:begin  
        addra4<=addra4+1;
	      k<=8'd97;
	     end
      8'd97:begin 
        if(i5<9)
	      begin 
	      i5<=i5+1;
	      k<=8'd95;
	      end
	      else
	      k<=8'd98;
	      end
      8'd98:begin 
         p2[j3]<=d[0]^d[1]^d[2]^d[3]^d[4]^d[5]^d[6]^d[7]^d[8]^d[9];
	      k<=8'd99;
	       end
	   8'd99:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd100;
		 end		 
	   8'd100:begin 
       if(j3<=9'd239) 
	    k<=8'd95;
	   else
	   begin
	   k<=8'd101;
	   end
	   end		
		8'd101:begin
        d[i5]<=bp2[douta4];
	     k<=8'd102;
	      end	
      8'd102:begin  
        addra4<=addra4+1;
	      k<=8'd103;
	     end
      8'd103:begin 
        if(i5<10)
	      begin 
	      i5<=i5+1;
	      k<=8'd101;
	      end
	      else
	      k<=8'd104;
	      end	  
      8'd104:begin 
         p2[j3]<=d[0]^d[1]^d[2]^d[3]^d[4]^d[5]^d[6]^d[7]^d[8]^d[9]^d[10];
	      k<=8'd105;
	       end
	   8'd105:begin 
	    j3<=j3+1;
		 i5<=4'd0;
		 k<=8'd106;
		 end
	   8'd106:begin 
       if(j3<=9'd263) 
	    k<=8'd101;
	   else
	   begin
	   k<=8'd107;
	   end
	   end
		8'd107:begin
		      u1<={p2,p1,u};
				k<=8'd108;
				end
		8'd108:begin 
		       out<=u1[j4];
				 k<=8'd109;
				 end
		8'd109:begin 
		       if(j4<575)
				 begin
				   j4<=j4+1;
					k<=8'd108;
					end
				 else
				   k<=8'd110;
					end
		default:k<=8'd110;				
	endcase
endmodule
