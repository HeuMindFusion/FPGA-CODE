`timescale 1ns / 1ps

module mux_10(
    input clk,
	 input rst,
	 input[7:0] mr,
	 input[7:0] r_9,
	 output[7:0] r_10
    );
wire[7:0] a_10;
reg[7:0] g_10;
reg[7:0] r10;

assign a_10 = mr;

 always @(posedge clk)                            //g10��m+r��ֵ���
  begin
  if(!rst)
   begin
	g_10<=0;
	r10<=0;
	end
  else
   begin
    g_10[0]<=a_10[2]^a_10[3]^a_10[4]^a_10[5]^a_10[6];	
	 g_10[1]<=a_10[0]^a_10[3]^a_10[4]^a_10[5]^a_10[6];	
	 g_10[2]<=a_10[0]^a_10[1]^a_10[2]^a_10[3]^a_10[6];	
    g_10[3]<=a_10[0]^a_10[1]^a_10[4]^a_10[5]^a_10[7];	
    g_10[4]<=a_10[0]^a_10[1]^a_10[3]^a_10[4]^a_10[5]^a_10[6]^a_10[7];	
	 g_10[5]<=a_10[0]^a_10[1]^a_10[2]^a_10[4]^a_10[5]^a_10[6]^a_10[7];	
	 g_10[6]<=a_10[0]^a_10[1]^a_10[2]^a_10[3]^a_10[5]^a_10[6]^a_10[7];	
	 g_10[7]<=a_10[1]^a_10[2]^a_10[3]^a_10[4]^a_10[6]^a_10[7];
	 r10<=r_9^g_10;
	end
 end

assign 	 r_10=r10;

endmodule
